library verilog;
use verilog.vl_types.all;
entity portadora_vlg_vec_tst is
end portadora_vlg_vec_tst;
